** sch_path: /usr/local/share/pdk/sky130A/libs.tech/xschem/sky130_tests/simulate_ff.sch
**.subckt simulate_ff CLEAR_ CLK
*.ipin CLEAR_
*.ipin CLK
x28 B[3] net4 net3 VGND VNB VPB VPWR net5 BNEXT[3] sky130_fd_sc_hd__fa_1
x33 B[2] net4 net2 VGND VNB VPB VPWR net3 BNEXT[2] sky130_fd_sc_hd__fa_1
x34 B[1] net4 net1 VGND VNB VPB VPWR net2 BNEXT[1] sky130_fd_sc_hd__fa_1
x35 B[0] CLEAR_ net4 VGND VNB VPB VPWR net1 BNEXT[0] sky130_fd_sc_hd__fa_1
x36 CLK net6 CLEAR_ VGND VNB VPB VPWR B[3] sky130_fd_sc_hd__dfrtp_1
x37 CLK net7 CLEAR_ VGND VNB VPB VPWR B[2] sky130_fd_sc_hd__dfrtp_1
x53 CLK net8 CLEAR_ VGND VNB VPB VPWR B[1] sky130_fd_sc_hd__dfrtp_1
x54 CLK net9 CLEAR_ VGND VNB VPB VPWR B[0] sky130_fd_sc_hd__dfrtp_1
x55 CLEAR_ VGND VNB VPB VPWR net4 sky130_fd_sc_hd__inv_2
x59 BNEXT[3] net10 VGND VNB VPB VPWR net6 sky130_fd_sc_hd__and2_1
x60 BNEXT[2] net10 VGND VNB VPB VPWR net7 sky130_fd_sc_hd__and2_1
x61 BNEXT[1] net10 VGND VNB VPB VPWR net8 sky130_fd_sc_hd__and2_1
x62 BNEXT[0] net10 VGND VNB VPB VPWR net9 sky130_fd_sc_hd__and2_1
x1 net10 VGND VNB VPB VPWR R sky130_fd_sc_hd__inv_2
x22 B[3] VGND VNB VPB VPWR net11 sky130_fd_sc_hd__inv_2
x23 B[2] VGND VNB VPB VPWR net12 sky130_fd_sc_hd__inv_2
x24 B[1] VGND VNB VPB VPWR net14 sky130_fd_sc_hd__inv_2
x25 B[0] VGND VNB VPB VPWR net13 sky130_fd_sc_hd__inv_2
x21 net11 net12 B[1] net13 VGND VNB VPB VPWR S[5] sky130_fd_sc_hd__nand4_1
x38 net17 net18 net19 net20 VGND VNB VPB VPWR S[1] sky130_fd_sc_hd__and4_1
x39 net11 net12 net14 B[0] VGND VNB VPB VPWR net15 sky130_fd_sc_hd__nand4_1
x40 net11 B[2] net14 net13 VGND VNB VPB VPWR net16 sky130_fd_sc_hd__nand4_1
x41 net15 net16 VGND VNB VPB VPWR S[0] sky130_fd_sc_hd__and2_1
x42 net11 net12 B[1] net13 VGND VNB VPB VPWR net18 sky130_fd_sc_hd__nand4_1
x43 net11 net12 B[1] B[0] VGND VNB VPB VPWR net19 sky130_fd_sc_hd__nand4_1
x44 net11 B[2] B[1] B[0] VGND VNB VPB VPWR net20 sky130_fd_sc_hd__nand4_1
x45 net11 net12 net14 B[0] VGND VNB VPB VPWR net17 sky130_fd_sc_hd__nand4_1
x46 net11 B[2] net14 B[0] VGND VNB VPB VPWR net21 sky130_fd_sc_hd__nand4_1
x47 net11 B[2] B[1] net13 VGND VNB VPB VPWR net22 sky130_fd_sc_hd__nand4_1
x48 net21 net22 VGND VNB VPB VPWR S[2] sky130_fd_sc_hd__and2_1
x49 net11 net12 net14 net13 VGND VNB VPB VPWR net23 sky130_fd_sc_hd__nand4_1
x50 net11 net12 net14 B[0] VGND VNB VPB VPWR net24 sky130_fd_sc_hd__nand4_1
x51 net11 B[2] B[1] B[0] VGND VNB VPB VPWR net25 sky130_fd_sc_hd__nand4_1
x52 net23 net24 net25 VGND VNB VPB VPWR S[3] sky130_fd_sc_hd__and3_1
x18 net11 net12 net14 net13 VGND VNB VPB VPWR net26 sky130_fd_sc_hd__and4_1
x19 net11 net12 B[1] net13 VGND VNB VPB VPWR net27 sky130_fd_sc_hd__and4_1
x20 net11 B[2] B[1] net13 VGND VNB VPB VPWR net28 sky130_fd_sc_hd__and4_1
x26 B[3] net12 net14 net13 VGND VNB VPB VPWR net29 sky130_fd_sc_hd__and4_1
x27 net26 net27 net28 net29 VGND VNB VPB VPWR S[4] sky130_fd_sc_hd__or4_1
x29 net11 net12 net14 B[0] VGND VNB VPB VPWR net30 sky130_fd_sc_hd__nand4_1
x30 net11 B[2] net14 net13 VGND VNB VPB VPWR net31 sky130_fd_sc_hd__nand4_1
x31 net11 B[2] B[1] B[0] VGND VNB VPB VPWR net32 sky130_fd_sc_hd__nand4_1
x32 net30 net31 net32 VGND VNB VPB VPWR S[6] sky130_fd_sc_hd__and3_1
x3 BNEXT[1] BNEXT[3] VGND VNB VPB VPWR net10 sky130_fd_sc_hd__nand2_1
**.ends
.end
