** sch_path: /home/oe23ranan/mpw/saradcspr2022/test.sch
**.subckt test
XR1 GND VDD GND sky130_fd_pr__res_high_po W=1 L=1 mult=1 m=1
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
