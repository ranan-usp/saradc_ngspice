** sch_path: /usr/local/share/pdk/sky130A/libs.tech/xschem/sky130_tests/test_stdcells.sch
**.subckt test_stdcells
x1 A B VSS VSS VCC VCC X sky130_fd_sc_hd__nand2_1
V1 A 0 pulse 0 1.8 '0.495/ 0.09e9 ' '0.01/0.09e9 ' '0.01/0.09e9 ' '0.49/0.09e9 ' '1/0.09e9 '
V2 B 0 pulse 0 1.8 '0.495/ 0.02e9 ' '0.01/0.02e9 ' '0.01/0.02e9 ' '0.49/0.02e9 ' '1/0.02e9 '
C1 X 0 3f m=1
x2 CLK A RESET_B VSS VSS VCC VCC Q sky130_fd_sc_hd__dfrtp_1
V3 CLK 0 pulse 0 1.8 '0.495/ 0.2e9 ' '0.01/0.2e9 ' '0.01/0.2e9 ' '0.49/0.2e9 ' '1/0.2e9 '
V4 RESET_B 0 pulse 0 1.8 '0.495/ 0.7e8 ' '0.01/0.7e8 ' '0.01/0.7e8 ' '0.49/0.7e8 ' '1/0.7e8 '
C2 Q 0 3f m=1
C3 Y 0 3f m=1
x3 A B VSS VSS VCC VCC Y sky130_fd_sc_hd__nor2b_1
x4 A CLK RESET_B VSS VSS VCC VCC Qlatch net1 sky130_fd_sc_hd__dlrbn_1
C4 Qlatch 0 3f m=1
x5 Y B VSS VSS VCC VCC net2 sky130_fd_sc_hd__nor2b_1
x6 net2 Qlatch VSS VSS VCC VCC net4 sky130_fd_sc_hd__nand2_1
x7 net3 net4 Q RESET_B VSS VSS VCC VCC XSCHEM sky130_fd_sc_hd__a31o_2
x8 Y VSS VSS VCC VCC net3 sky130_fd_sc_hd__inv_2
**** begin user architecture code


.options acct list
.temp 25
vvcc vcc 0 dc 1.8
vvss vss 0 0
.control
tran 30p 80n
plot a b+2 clk+4 reset_b+6 x+8 y+10 q+12 qlatch+14
write test_stdcells.raw
.endc


 .lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
**.ends
.end
